LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;

-- GRUPO:
-- Bruno Pereira Bannwart
-- Luis Marcelo Stein d'Avila

ENTITY CPU IS
	PORT (
		Clock, Resetn	:IN	STD_LOGIC
	);
END CPU;

ARCHITECTURE Behavior OF CPU IS 

	
	
	--PC
	SIGNAL Address: STD_LOGIC_VECTOR(15 DOWNTO 0);
	
	--CACHE
	SIGNAL instruction	:	STD_LOGIC_VECTOR(15 DOWNTO 0);
	
	-- IF_ID
	SIGNAL Ime			:  STD_LOGIC;
	SIGNAL OPcode		:  STD_LOGIC_vECTOR(2 DOWNTO 0);
	SIGNAL Ri			:	STD_LOGIC_vECTOR(3 DOWNTO 0);
	SIGNAL Rj			:	STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL Rk_ime		:	STD_LOGIC_VECTOR(3 DOWNTO 0);
	
	--Unidade de Controle
	SIGNAL UCOUT : STD_LOGIC_VECTOR (3 DOWNTO 0);
	
	--ID_EX
	
	SIGNAL Q1	: STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL Q2	: STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL WB	: STD_LOGIC_VECTOR(4 DOWNTO 0);
	SIGNAL ALUOp :  STD_LOGIC_VECTOR(1 DOWNTO 0);
	SIGNAL Cin :  STD_LOGIC;
	
	
	--RegBank
	SIGNAL RegA	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL RegB	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	
	--MUX2
	SIGNAL Operator2 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	
	--ULA
	SIGNAL Result		:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL Overflow	:	STD_LOGIC;
	SIGNAL Cout 		:	STD_LOGIC;
	
	--EX_WB
	
	SIGNAL WBResult	: STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL RegDst: STD_LOGIC_VECTOR (3 DOWNTO 0);
	SIGNAL Regwrite:  STD_LOGIC;
	
	-- Todos os componentes necessarios da ula
	
	COMPONENT PC
		PORT (
			Address_out				 : 	OUT 	STD_LOGIC_VECTOR(15 DOWNTO 0);
			Clock,Resetn : 	IN 	STD_LOGIC
		);
	END COMPONENT PC;
	
	COMPONENT RegBank
		PORT (
			regwrite, Clock, Resetn: IN STD_LOGIC;
			S1: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
			S2: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
			N: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
			Rs: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			Rt: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			Rd: IN STD_LOGIC_VECTOR (3 DOWNTO 0)
		);
	END COMPONENT RegBank;	
	
	COMPONENT ULA
		PORT (
			Cin, Clock  	:	IN  STD_LOGIC;
			X,Y  				:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
			S    				:	OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			Op   				:	IN STD_LOGIC_VECTOR(1 DOWNTO 0);
			Cout,Overflow 	: 	OUT STD_LOGIC
		);
	END COMPONENT ULA;
	
	COMPONENT CACHE
	PORT (
		address_PC: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		data_instruction :OUT STD_LOGIC_VECTOR (15 DOWNTO 0); 
		Clock: IN STD_LOGIC
	);
	END COMPONENT CACHE;
	
	COMPONENT MUX_EXT
		PORT(
		X: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		Y: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		Z: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
		S, Clock: STD_LOGIC
	);
	END COMPONENT MUX_EXT;
	
	COMPONENT Controle IS
	PORT (
		instruction		:IN 	STD_LOGIC_VECTOR(2 DOWNTO 0);
		Resetn, Clock		:IN STD_LOGIC;
		UCOut: OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
		
	);
	END COMPONENT Controle;

	COMPONENT IF_ID
		PORT (
		Mem_in: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		Resetn: IN STD_LOGIC;
			Ri, Rj, Rk: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
			OpCode: OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
			Ime: OUT STD_LOGIC;
			Clock: IN STD_LOGIC
			);
	END COMPONENT IF_ID;
	
	COMPONENT ID_EX
	PORT (
			D1	:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			D2	:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			UC :IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			RegDst :IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			Resetn, Clock :IN STD_LOGIC;
			Q1	:OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			Q2	:OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			WB	:OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
			ALUOp : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
			Cin : OUT STD_LOGIC
			
			);
	END COMPONENT ID_EX;
	
	COMPONENT EX_WB
	PORT (
			D	:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			Resetn, Clock :IN STD_LOGIC;
			WB	:IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			Q1	:OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			RegDst: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
			Regwrite: OUT STD_LOGIC
			
			);
	END COMPONENT EX_WB;
	
BEGIN
	PC1:  PC PORT MAP(Address, Clock, Resetn);
	
	CACHE1: CACHE PORT MAP(Address, instruction, Clock);
	
	IF_ID1: IF_ID PORT MAP(Instruction, Resetn, Ri, Rj, Rk_ime, OPcode, Ime, Clock);
	
	UC1: Controle PORT MAP(OPCode, Resetn, Clock, UCOut); 
	
	RB: RegBank PORT MAP(RegWrite, Clock, Resetn, RegA, RegB, WBResult, Rj, Rk_ime, RegDst);
	
	MUX1: MUX_EXT PORT MAP (RegB, Rk_ime, Operator2, Ime, Clock);
	
	ID_EX1: ID_EX PORT MAP (RegA, Operator2, UCOut,Ri, Resetn, Clock, Q1, Q2, WB, ALUOp, Cin); --alterar aqui
	
	ULA1 : ULA PORT MAP (Cin, Clock, Q1, Q2, Result, ALUOp, Cout, Overflow);
	
	EX_WB1: EX_WB PORT MAP (Result, Resetn, Clock, WB, WBResult,RegDst, RegWrite);
	
	END Behavior;
		
	